module displaytest(wei,duan);
output wei;
output duan;

endmodule
