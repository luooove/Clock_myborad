module displaytest(Wei,Duan);
output[7:0] Wei;
output[7:0] Duan;

assign Duan = 8'b1101_1010;
assign Wei = 8'b0000_0000;


endmodule
